-- megafunction wizard: %ALTMEMMULT%
-- GENERATION: STANDARD
-- VERSION: WM1.0
-- MODULE: altmemmult 

-- ============================================================
-- File Name: memmult.vhd
-- Megafunction Name(s):
-- 			altmemmult
--
-- Simulation Library Files(s):
-- 			altera_mf;cyclone
-- ============================================================
-- ************************************************************
-- THIS IS A WIZARD-GENERATED FILE. DO NOT EDIT THIS FILE!
--
-- 7.1 Build 156 04/30/2007 SJ Web Edition
-- ************************************************************


--Copyright (C) 1991-2007 Altera Corporation
--Your use of Altera Corporation's design tools, logic functions 
--and other software and tools, and its AMPP partner logic 
--functions, and any output files from any of the foregoing 
--(including device programming or simulation files), and any 
--associated documentation or information are expressly subject 
--to the terms and conditions of the Altera Program License 
--Subscription Agreement, Altera MegaCore Function License 
--Agreement, or other applicable license agreement, including, 
--without limitation, that your use is for the sole purpose of 
--programming logic devices manufactured by Altera and sold by 
--Altera or its authorized distributors.  Please refer to the 
--applicable agreement for further details.


--altmemmult CBX_AUTO_BLACKBOX="ALL" COEFF_REPRESENTATION="SIGNED" COEFFICIENT0="1234" DATA_REPRESENTATION="SIGNED" DEVICE_FAMILY="Cyclone" MAX_CLOCK_CYCLES_PER_RESULT=8 RAM_BLOCK_TYPE="AUTO" TOTAL_LATENCY=11 WIDTH_C=32 WIDTH_D=32 WIDTH_R=64 clock data_in result result_valid sload_data
--VERSION_BEGIN 7.1 cbx_altaccumulate 2006:05:24:11:25:36:SJ cbx_altmemmult 2007:01:23:15:28:00:SJ cbx_altsyncram 2007:03:22:08:29:24:SJ cbx_cycloneii 2007:01:23:09:39:40:SJ cbx_lpm_add_sub 2007:01:08:11:15:18:SJ cbx_lpm_compare 2007:02:05:11:33:54:SJ cbx_lpm_counter 2007:03:22:23:17:10:SJ cbx_lpm_decode 2006:11:21:10:27:00:SJ cbx_lpm_mux 2006:11:21:10:27:10:SJ cbx_mgl 2007:04:03:14:06:46:SJ cbx_stratix 2007:04:12:16:43:52:SJ cbx_stratixii 2007:02:12:17:08:26:SJ cbx_stratixiii 2007:03:13:14:47:12:SJ cbx_util_mgl 2007:01:15:12:22:48:SJ  VERSION_END


--alt_abs CBX_AUTO_BLACKBOX="ALL" DEVICE_FAMILY="Cyclone" LPM_WIDTH=4 abs clock data result sign_bit sload sload_data
--VERSION_BEGIN 7.1 cbx_altaccumulate 2006:05:24:11:25:36:SJ cbx_altmemmult 2007:01:23:15:28:00:SJ cbx_altsyncram 2007:03:22:08:29:24:SJ cbx_cycloneii 2007:01:23:09:39:40:SJ cbx_lpm_add_sub 2007:01:08:11:15:18:SJ cbx_lpm_compare 2007:02:05:11:33:54:SJ cbx_lpm_counter 2007:03:22:23:17:10:SJ cbx_lpm_decode 2006:11:21:10:27:00:SJ cbx_lpm_mux 2006:11:21:10:27:10:SJ cbx_mgl 2007:04:03:14:06:46:SJ cbx_stratix 2007:04:12:16:43:52:SJ cbx_stratixii 2007:02:12:17:08:26:SJ cbx_stratixiii 2007:03:13:14:47:12:SJ cbx_util_mgl 2007:01:15:12:22:48:SJ  VERSION_END

 LIBRARY cyclone;
 USE cyclone.all;

--synthesis_resources = lut 5 
 LIBRARY ieee;
 USE ieee.std_logic_1164.all;

 ENTITY  memmult_abs_bla IS 
	 PORT 
	 ( 
		 a_abs	:	IN  STD_LOGIC;
		 clock	:	IN  STD_LOGIC;
		 data	:	IN  STD_LOGIC_VECTOR (3 DOWNTO 0);
		 result	:	OUT  STD_LOGIC_VECTOR (3 DOWNTO 0);
		 sign_bit	:	IN  STD_LOGIC := '0';
		 sload	:	IN  STD_LOGIC := '0';
		 sload_data	:	IN  STD_LOGIC_VECTOR (3 DOWNTO 0)
	 ); 
 END memmult_abs_bla;

 ARCHITECTURE RTL OF memmult_abs_bla IS

	 ATTRIBUTE synthesis_clearbox : boolean;
	 ATTRIBUTE synthesis_clearbox OF RTL : ARCHITECTURE IS true;
	 SIGNAL	 inv_reg	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL  wire_strx_lcell9a_0cout	:	STD_LOGIC;
	 SIGNAL  wire_strx_lcell9a_1cout	:	STD_LOGIC;
	 SIGNAL  wire_strx_lcell9a_2cout	:	STD_LOGIC;
	 SIGNAL  wire_strx_lcell9a_dataa	:	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  wire_strx_lcell9a_datab	:	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  wire_strx_lcell9a_datac	:	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  wire_strx_lcell9a_regout	:	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 COMPONENT  cyclone_lcell
	 GENERIC 
	 (
		cin0_used	:	STRING := "false";
		cin1_used	:	STRING := "false";
		cin_used	:	STRING := "false";
		lut_mask	:	STRING;
		operation_mode	:	STRING := "normal";
		output_mode	:	STRING := "reg_and_comb";
		power_up	:	STRING := "low";
		register_cascade_mode	:	STRING := "off";
		sum_lutc_input	:	STRING := "datac";
		synch_mode	:	STRING := "off";
		x_on_violation	:	STRING := "on";
		lpm_type	:	STRING := "cyclone_lcell"
	 );
	 PORT
	 ( 
		aclr	:	IN STD_LOGIC := '0';
		aload	:	IN STD_LOGIC := '0';
		cin	:	IN STD_LOGIC := '0';
		clk	:	IN STD_LOGIC := '0';
		combout	:	OUT STD_LOGIC;
		cout	:	OUT STD_LOGIC;
		dataa	:	IN STD_LOGIC := '1';
		datab	:	IN STD_LOGIC := '1';
		datac	:	IN STD_LOGIC := '1';
		datad	:	IN STD_LOGIC := '1';
		ena	:	IN STD_LOGIC := '1';
		inverta	:	IN STD_LOGIC := '0';
		regcascin	:	IN STD_LOGIC := '0';
		regout	:	OUT STD_LOGIC;
		sclr	:	IN STD_LOGIC := '0';
		sload	:	IN STD_LOGIC := '0'
	 ); 
	 END COMPONENT;
 BEGIN

	result <= wire_strx_lcell9a_regout;
	PROCESS (clock)
	BEGIN
		IF (clock = '1' AND clock'event) THEN inv_reg <= (a_abs AND sign_bit);
		END IF;
	END PROCESS;
	wire_strx_lcell9a_dataa <= data;
	wire_strx_lcell9a_datab <= "0000";
	wire_strx_lcell9a_datac <= sload_data;
	strx_lcell9a_0 :  cyclone_lcell
	  GENERIC MAP (
		cin_used => "false",
		lut_mask => "96E8",
		operation_mode => "arithmetic",
		sum_lutc_input => "cin",
		synch_mode => "on"
	  )
	  PORT MAP ( 
		clk => clock,
		cout => wire_strx_lcell9a_0cout,
		dataa => wire_strx_lcell9a_dataa(0),
		datab => wire_strx_lcell9a_datab(0),
		datac => wire_strx_lcell9a_datac(0),
		inverta => inv_reg,
		regout => wire_strx_lcell9a_regout(0),
		sload => sload
	  );
	strx_lcell9a_1 :  cyclone_lcell
	  GENERIC MAP (
		cin_used => "true",
		lut_mask => "96E8",
		operation_mode => "arithmetic",
		sum_lutc_input => "cin",
		synch_mode => "on"
	  )
	  PORT MAP ( 
		cin => wire_strx_lcell9a_0cout,
		clk => clock,
		cout => wire_strx_lcell9a_1cout,
		dataa => wire_strx_lcell9a_dataa(1),
		datab => wire_strx_lcell9a_datab(1),
		datac => wire_strx_lcell9a_datac(1),
		inverta => inv_reg,
		regout => wire_strx_lcell9a_regout(1),
		sload => sload
	  );
	strx_lcell9a_2 :  cyclone_lcell
	  GENERIC MAP (
		cin_used => "true",
		lut_mask => "96E8",
		operation_mode => "arithmetic",
		sum_lutc_input => "cin",
		synch_mode => "on"
	  )
	  PORT MAP ( 
		cin => wire_strx_lcell9a_1cout,
		clk => clock,
		cout => wire_strx_lcell9a_2cout,
		dataa => wire_strx_lcell9a_dataa(2),
		datab => wire_strx_lcell9a_datab(2),
		datac => wire_strx_lcell9a_datac(2),
		inverta => inv_reg,
		regout => wire_strx_lcell9a_regout(2),
		sload => sload
	  );
	strx_lcell9a_3 :  cyclone_lcell
	  GENERIC MAP (
		cin_used => "true",
		lut_mask => "9696",
		operation_mode => "normal",
		sum_lutc_input => "cin",
		synch_mode => "on"
	  )
	  PORT MAP ( 
		cin => wire_strx_lcell9a_2cout,
		clk => clock,
		dataa => wire_strx_lcell9a_dataa(3),
		datab => wire_strx_lcell9a_datab(3),
		datac => wire_strx_lcell9a_datac(3),
		inverta => inv_reg,
		regout => wire_strx_lcell9a_regout(3),
		sload => sload
	  );

 END RTL; --memmult_abs_bla


--altshiftreg CBX_AUTO_BLACKBOX="ALL" LPM_DIRECTION="RIGHT" LPM_WIDTH=28 SHIFT_DISTANCE=4 clock data load shiftout
--VERSION_BEGIN 7.1 cbx_altaccumulate 2006:05:24:11:25:36:SJ cbx_altmemmult 2007:01:23:15:28:00:SJ cbx_altsyncram 2007:03:22:08:29:24:SJ cbx_cycloneii 2007:01:23:09:39:40:SJ cbx_lpm_add_sub 2007:01:08:11:15:18:SJ cbx_lpm_compare 2007:02:05:11:33:54:SJ cbx_lpm_counter 2007:03:22:23:17:10:SJ cbx_lpm_decode 2006:11:21:10:27:00:SJ cbx_lpm_mux 2006:11:21:10:27:10:SJ cbx_mgl 2007:04:03:14:06:46:SJ cbx_stratix 2007:04:12:16:43:52:SJ cbx_stratixii 2007:02:12:17:08:26:SJ cbx_stratixiii 2007:03:13:14:47:12:SJ cbx_util_mgl 2007:01:15:12:22:48:SJ  VERSION_END

--synthesis_resources = lut 28 
 LIBRARY ieee;
 USE ieee.std_logic_1164.all;

 ENTITY  memmult_altshiftreg_tda IS 
	 PORT 
	 ( 
		 clock	:	IN  STD_LOGIC;
		 data	:	IN  STD_LOGIC_VECTOR (27 DOWNTO 0) := (OTHERS => '0');
		 load	:	IN  STD_LOGIC := '0';
		 q	:	OUT  STD_LOGIC_VECTOR (27 DOWNTO 0);
		 shiftout	:	OUT  STD_LOGIC_VECTOR (3 DOWNTO 0)
	 ); 
 END memmult_altshiftreg_tda;

 ARCHITECTURE RTL OF memmult_altshiftreg_tda IS

	 ATTRIBUTE synthesis_clearbox : boolean;
	 ATTRIBUTE synthesis_clearbox OF RTL : ARCHITECTURE IS true;
	 SIGNAL	 dffe10a	:	STD_LOGIC_VECTOR(27 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL  wire_altshiftreg1_w_lg_w_lg_load70w71w	:	STD_LOGIC_VECTOR (27 DOWNTO 0);
	 SIGNAL  wire_altshiftreg1_w_lg_w_lg_sclr74w75w	:	STD_LOGIC_VECTOR (27 DOWNTO 0);
	 SIGNAL  wire_altshiftreg1_w_lg_load69w	:	STD_LOGIC_VECTOR (27 DOWNTO 0);
	 SIGNAL  wire_altshiftreg1_w_lg_load70w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altshiftreg1_w_lg_sclr74w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altshiftreg1_w_lg_w_lg_w_lg_load70w71w72w	:	STD_LOGIC_VECTOR (27 DOWNTO 0);
	 SIGNAL  wire_altshiftreg1_w_lg_sset73w	:	STD_LOGIC_VECTOR (27 DOWNTO 0);
	 SIGNAL  sclr	:	STD_LOGIC;
	 SIGNAL  shift_node :	STD_LOGIC_VECTOR (27 DOWNTO 0);
	 SIGNAL  shiftin_wire :	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  sset	:	STD_LOGIC;
 BEGIN

	loop0 : FOR i IN 0 TO 27 GENERATE 
		wire_altshiftreg1_w_lg_w_lg_load70w71w(i) <= wire_altshiftreg1_w_lg_load70w(0) AND shift_node(i);
	END GENERATE loop0;
	loop1 : FOR i IN 0 TO 27 GENERATE 
		wire_altshiftreg1_w_lg_w_lg_sclr74w75w(i) <= wire_altshiftreg1_w_lg_sclr74w(0) AND wire_altshiftreg1_w_lg_sset73w(i);
	END GENERATE loop1;
	loop2 : FOR i IN 0 TO 27 GENERATE 
		wire_altshiftreg1_w_lg_load69w(i) <= load AND data(i);
	END GENERATE loop2;
	wire_altshiftreg1_w_lg_load70w(0) <= NOT load;
	wire_altshiftreg1_w_lg_sclr74w(0) <= NOT sclr;
	loop3 : FOR i IN 0 TO 27 GENERATE 
		wire_altshiftreg1_w_lg_w_lg_w_lg_load70w71w72w(i) <= wire_altshiftreg1_w_lg_w_lg_load70w71w(i) OR wire_altshiftreg1_w_lg_load69w(i);
	END GENERATE loop3;
	loop4 : FOR i IN 0 TO 27 GENERATE 
		wire_altshiftreg1_w_lg_sset73w(i) <= sset OR wire_altshiftreg1_w_lg_w_lg_w_lg_load70w71w72w(i);
	END GENERATE loop4;
	q <= dffe10a;
	sclr <= '0';
	shift_node <= ( shiftin_wire & dffe10a(27 DOWNTO 4));
	shiftin_wire <= "0000";
	shiftout <= dffe10a(3 DOWNTO 0);
	sset <= '0';
	PROCESS (clock)
	BEGIN
		IF (clock = '1' AND clock'event) THEN dffe10a <= wire_altshiftreg1_w_lg_w_lg_sclr74w75w;
		END IF;
	END PROCESS;

 END RTL; --memmult_altshiftreg_tda


--altshiftreg CBX_AUTO_BLACKBOX="ALL" LPM_DIRECTION="RIGHT" LPM_WIDTH=28 SHIFT_DISTANCE=4 clock q shiftin
--VERSION_BEGIN 7.1 cbx_altaccumulate 2006:05:24:11:25:36:SJ cbx_altmemmult 2007:01:23:15:28:00:SJ cbx_altsyncram 2007:03:22:08:29:24:SJ cbx_cycloneii 2007:01:23:09:39:40:SJ cbx_lpm_add_sub 2007:01:08:11:15:18:SJ cbx_lpm_compare 2007:02:05:11:33:54:SJ cbx_lpm_counter 2007:03:22:23:17:10:SJ cbx_lpm_decode 2006:11:21:10:27:00:SJ cbx_lpm_mux 2006:11:21:10:27:10:SJ cbx_mgl 2007:04:03:14:06:46:SJ cbx_stratix 2007:04:12:16:43:52:SJ cbx_stratixii 2007:02:12:17:08:26:SJ cbx_stratixiii 2007:03:13:14:47:12:SJ cbx_util_mgl 2007:01:15:12:22:48:SJ  VERSION_END

--synthesis_resources = lut 28 
 LIBRARY ieee;
 USE ieee.std_logic_1164.all;

 ENTITY  memmult_altshiftreg_ji9 IS 
	 PORT 
	 ( 
		 clock	:	IN  STD_LOGIC;
		 q	:	OUT  STD_LOGIC_VECTOR (27 DOWNTO 0);
		 shiftin	:	IN  STD_LOGIC_VECTOR (3 DOWNTO 0) := (OTHERS => '1');
		 shiftout	:	OUT  STD_LOGIC_VECTOR (3 DOWNTO 0)
	 ); 
 END memmult_altshiftreg_ji9;

 ARCHITECTURE RTL OF memmult_altshiftreg_ji9 IS

	 ATTRIBUTE synthesis_clearbox : boolean;
	 ATTRIBUTE synthesis_clearbox OF RTL : ARCHITECTURE IS true;
	 SIGNAL	 dffe11a	:	STD_LOGIC_VECTOR(27 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL  wire_altshiftreg8_w_lg_w_lg_load80w81w	:	STD_LOGIC_VECTOR (27 DOWNTO 0);
	 SIGNAL  wire_altshiftreg8_w_lg_w_lg_sclr84w85w	:	STD_LOGIC_VECTOR (27 DOWNTO 0);
	 SIGNAL  wire_altshiftreg8_w_lg_load79w	:	STD_LOGIC_VECTOR (27 DOWNTO 0);
	 SIGNAL  wire_altshiftreg8_w_lg_load80w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altshiftreg8_w_lg_sclr84w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altshiftreg8_w_lg_w_lg_w_lg_load80w81w82w	:	STD_LOGIC_VECTOR (27 DOWNTO 0);
	 SIGNAL  wire_altshiftreg8_w_lg_sset83w	:	STD_LOGIC_VECTOR (27 DOWNTO 0);
	 SIGNAL  data	:	STD_LOGIC_VECTOR (27 DOWNTO 0);
	 SIGNAL  load	:	STD_LOGIC;
	 SIGNAL  sclr	:	STD_LOGIC;
	 SIGNAL  shift_node :	STD_LOGIC_VECTOR (27 DOWNTO 0);
	 SIGNAL  shiftin_wire :	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  sset	:	STD_LOGIC;
 BEGIN

	loop5 : FOR i IN 0 TO 27 GENERATE 
		wire_altshiftreg8_w_lg_w_lg_load80w81w(i) <= wire_altshiftreg8_w_lg_load80w(0) AND shift_node(i);
	END GENERATE loop5;
	loop6 : FOR i IN 0 TO 27 GENERATE 
		wire_altshiftreg8_w_lg_w_lg_sclr84w85w(i) <= wire_altshiftreg8_w_lg_sclr84w(0) AND wire_altshiftreg8_w_lg_sset83w(i);
	END GENERATE loop6;
	loop7 : FOR i IN 0 TO 27 GENERATE 
		wire_altshiftreg8_w_lg_load79w(i) <= load AND data(i);
	END GENERATE loop7;
	wire_altshiftreg8_w_lg_load80w(0) <= NOT load;
	wire_altshiftreg8_w_lg_sclr84w(0) <= NOT sclr;
	loop8 : FOR i IN 0 TO 27 GENERATE 
		wire_altshiftreg8_w_lg_w_lg_w_lg_load80w81w82w(i) <= wire_altshiftreg8_w_lg_w_lg_load80w81w(i) OR wire_altshiftreg8_w_lg_load79w(i);
	END GENERATE loop8;
	loop9 : FOR i IN 0 TO 27 GENERATE 
		wire_altshiftreg8_w_lg_sset83w(i) <= sset OR wire_altshiftreg8_w_lg_w_lg_w_lg_load80w81w82w(i);
	END GENERATE loop9;
	data <= (OTHERS => '0');
	load <= '0';
	q <= dffe11a;
	sclr <= '0';
	shift_node <= ( shiftin_wire & dffe11a(27 DOWNTO 4));
	shiftin_wire <= shiftin;
	shiftout <= dffe11a(3 DOWNTO 0);
	sset <= '0';
	PROCESS (clock)
	BEGIN
		IF (clock = '1' AND clock'event) THEN dffe11a <= wire_altshiftreg8_w_lg_w_lg_sclr84w85w;
		END IF;
	END PROCESS;

 END RTL; --memmult_altshiftreg_ji9

 LIBRARY altera_mf;
 USE altera_mf.all;

--synthesis_resources = altaccumulate 1 altsyncram 1 lut 82 
 LIBRARY ieee;
 USE ieee.std_logic_1164.all;

 ENTITY  memmult_altmemmult_v6q IS 
	 PORT 
	 ( 
		 clock	:	IN  STD_LOGIC;
		 data_in	:	IN  STD_LOGIC_VECTOR (31 DOWNTO 0);
		 result	:	OUT  STD_LOGIC_VECTOR (63 DOWNTO 0);
		 result_valid	:	OUT  STD_LOGIC;
		 sload_data	:	IN  STD_LOGIC := '0'
	 ); 
 END memmult_altmemmult_v6q;

 ARCHITECTURE RTL OF memmult_altmemmult_v6q IS

	 ATTRIBUTE synthesis_clearbox : boolean;
	 ATTRIBUTE synthesis_clearbox OF RTL : ARCHITECTURE IS true;
	 SIGNAL  wire_abs3_data	:	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  wire_abs3_result	:	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  wire_abs3_sign_bit	:	STD_LOGIC;
	 SIGNAL  wire_abs3_sload_data	:	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  wire_accum7_add_sub	:	STD_LOGIC;
	 SIGNAL  wire_dffe4a_w_lg_w_q_range54w55w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_accum7_data	:	STD_LOGIC_VECTOR (35 DOWNTO 0);
	 SIGNAL  wire_accum7_result	:	STD_LOGIC_VECTOR (36 DOWNTO 0);
	 SIGNAL  wire_altshiftreg1_data	:	STD_LOGIC_VECTOR (27 DOWNTO 0);
	 SIGNAL  wire_altshiftreg1_q	:	STD_LOGIC_VECTOR (27 DOWNTO 0);
	 SIGNAL  wire_altshiftreg1_shiftout	:	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  wire_altshiftreg8_q	:	STD_LOGIC_VECTOR (27 DOWNTO 0);
	 SIGNAL  wire_altshiftreg8_shiftout	:	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  wire_altsyncram6_q_a	:	STD_LOGIC_VECTOR (35 DOWNTO 0);
	 SIGNAL	 dffe2a0	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 dffe2a1	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 dffe2a2	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL  wire_dffe2a_w_lg_q9w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL	 dffe2a3	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL  wire_dffe2a_w_lg_q10w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL	 dffe2a4	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL  wire_dffe2a_w_lg_q12w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL	 dffe2a5	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL  wire_dffe2a_w_lg_q14w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL	 dffe2a6	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL  wire_dffe2a_w_lg_q16w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL	 dffe2a7	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL  wire_dffe2a_w_lg_q18w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL	 dffe2a8	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL  wire_dffe2a_w_lg_q20w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL	 dffe2a9	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL  wire_dffe2a_w_lg_q22w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL	 dffe2a10	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 dffe4a	:	STD_LOGIC_VECTOR(3 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL  wire_dffe4a_w44w	:	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL	 dffe5a0	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL  wire_dffe5a_w_lg_q32w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL	 dffe5a1	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL  wire_dffe5a_w_lg_q34w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL	 dffe5a2	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL  wire_dffe5a_w_lg_q36w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL	 dffe5a3	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL  wire_dffe5a_w_lg_q38w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL	 dffe5a4	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL  wire_dffe5a_w_lg_q40w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL	 dffe5a5	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL  wire_dffe5a_w_lg_q42w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_sclr4w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_sload_data31w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  result_wire :	STD_LOGIC_VECTOR (63 DOWNTO 0);
	 SIGNAL  sclr	:	STD_LOGIC;
	 COMPONENT  memmult_abs_bla
	 PORT
	 ( 
		a_abs	:	IN  STD_LOGIC;
		clock	:	IN  STD_LOGIC;
		data	:	IN  STD_LOGIC_VECTOR(3 DOWNTO 0);
		result	:	OUT  STD_LOGIC_VECTOR(3 DOWNTO 0);
		sign_bit	:	IN  STD_LOGIC := '0';
		sload	:	IN  STD_LOGIC := '0';
		sload_data	:	IN  STD_LOGIC_VECTOR(3 DOWNTO 0)
	 ); 
	 END COMPONENT;
	 COMPONENT  altaccumulate
	 GENERIC 
	 (
		CARRY_CHAIN	:	STRING := "MANUAL";
		CARRY_CHAIN_LENGTH	:	NATURAL := 32;
		EXTRA_LATENCY	:	NATURAL := 0;
		LPM_REPRESENTATION	:	STRING := "UNSIGNED";
		RIGHT_SHIFT_DISTANCE	:	NATURAL := 0;
		USE_WYS	:	STRING := "ON";
		WIDTH_IN	:	NATURAL;
		WIDTH_OUT	:	NATURAL;
		lpm_type	:	STRING := "altaccumulate"
	 );
	 PORT
	 ( 
		aclr	:	IN STD_LOGIC := '0';
		add_sub	:	IN STD_LOGIC := '1';
		cin	:	IN STD_LOGIC := 'Z';
		clken	:	IN STD_LOGIC := '1';
		clock	:	IN STD_LOGIC;
		cout	:	OUT STD_LOGIC;
		data	:	IN STD_LOGIC_VECTOR(WIDTH_IN-1 DOWNTO 0);
		overflow	:	OUT STD_LOGIC;
		result	:	OUT STD_LOGIC_VECTOR(WIDTH_OUT-1 DOWNTO 0);
		sign_data	:	IN STD_LOGIC := '0';
		sload	:	IN STD_LOGIC := '0'
	 ); 
	 END COMPONENT;
	 COMPONENT  memmult_altshiftreg_tda
	 PORT
	 ( 
		clock	:	IN  STD_LOGIC;
		data	:	IN  STD_LOGIC_VECTOR(27 DOWNTO 0) := (OTHERS => '0');
		load	:	IN  STD_LOGIC := '0';
		q	:	OUT  STD_LOGIC_VECTOR(27 DOWNTO 0);
		shiftout	:	OUT  STD_LOGIC_VECTOR(3 DOWNTO 0)
	 ); 
	 END COMPONENT;
	 COMPONENT  memmult_altshiftreg_ji9
	 PORT
	 ( 
		clock	:	IN  STD_LOGIC;
		q	:	OUT  STD_LOGIC_VECTOR(27 DOWNTO 0);
		shiftin	:	IN  STD_LOGIC_VECTOR(3 DOWNTO 0) := (OTHERS => '1');
		shiftout	:	OUT  STD_LOGIC_VECTOR(3 DOWNTO 0)
	 ); 
	 END COMPONENT;
	 COMPONENT  altsyncram
	 GENERIC 
	 (
		ADDRESS_ACLR_A	:	STRING := "UNUSED";
		ADDRESS_ACLR_B	:	STRING := "NONE";
		ADDRESS_REG_B	:	STRING := "CLOCK1";
		BYTE_SIZE	:	NATURAL := 8;
		BYTEENA_ACLR_A	:	STRING := "UNUSED";
		BYTEENA_ACLR_B	:	STRING := "NONE";
		BYTEENA_REG_B	:	STRING := "CLOCK1";
		CLOCK_ENABLE_CORE_A	:	STRING := "USE_INPUT_CLKEN";
		CLOCK_ENABLE_CORE_B	:	STRING := "USE_INPUT_CLKEN";
		CLOCK_ENABLE_INPUT_A	:	STRING := "NORMAL";
		CLOCK_ENABLE_INPUT_B	:	STRING := "NORMAL";
		CLOCK_ENABLE_OUTPUT_A	:	STRING := "NORMAL";
		CLOCK_ENABLE_OUTPUT_B	:	STRING := "NORMAL";
		ENABLE_ECC	:	STRING := "FALSE";
		IMPLEMENT_IN_LES	:	STRING := "OFF";
		INDATA_ACLR_A	:	STRING := "UNUSED";
		INDATA_ACLR_B	:	STRING := "NONE";
		INDATA_REG_B	:	STRING := "CLOCK1";
		INIT_FILE	:	STRING := "UNUSED";
		INIT_FILE_LAYOUT	:	STRING := "PORT_A";
		MAXIMUM_DEPTH	:	NATURAL := 0;
		NUMWORDS_A	:	NATURAL := 0;
		NUMWORDS_B	:	NATURAL := 0;
		OPERATION_MODE	:	STRING := "BIDIR_DUAL_PORT";
		OUTDATA_ACLR_A	:	STRING := "NONE";
		OUTDATA_ACLR_B	:	STRING := "NONE";
		OUTDATA_REG_A	:	STRING := "UNREGISTERED";
		OUTDATA_REG_B	:	STRING := "UNREGISTERED";
		POWER_UP_UNINITIALIZED	:	STRING := "FALSE";
		RAM_BLOCK_TYPE	:	STRING := "AUTO";
		RDCONTROL_ACLR_B	:	STRING := "NONE";
		RDCONTROL_REG_B	:	STRING := "CLOCK1";
		READ_DURING_WRITE_MODE_MIXED_PORTS	:	STRING := "DONT_CARE";
		read_during_write_mode_port_a	:	STRING := "NEW_DATA_NO_NBE_READ";
		read_during_write_mode_port_b	:	STRING := "NEW_DATA_NO_NBE_READ";
		WIDTH_A	:	NATURAL;
		WIDTH_B	:	NATURAL := 1;
		WIDTH_BYTEENA_A	:	NATURAL := 1;
		WIDTH_BYTEENA_B	:	NATURAL := 1;
		WIDTHAD_A	:	NATURAL;
		WIDTHAD_B	:	NATURAL := 1;
		WRCONTROL_ACLR_A	:	STRING := "UNUSED";
		WRCONTROL_ACLR_B	:	STRING := "NONE";
		WRCONTROL_WRADDRESS_REG_B	:	STRING := "CLOCK1";
		INTENDED_DEVICE_FAMILY	:	STRING := "Cyclone";
		lpm_hint	:	STRING := "UNUSED";
		lpm_type	:	STRING := "altsyncram"
	 );
	 PORT
	 ( 
		aclr0	:	IN STD_LOGIC := '0';
		aclr1	:	IN STD_LOGIC := '0';
		address_a	:	IN STD_LOGIC_VECTOR(WIDTHAD_A-1 DOWNTO 0);
		address_b	:	IN STD_LOGIC_VECTOR(WIDTHAD_B-1 DOWNTO 0) := (OTHERS => '1');
		addressstall_a	:	IN STD_LOGIC := '0';
		addressstall_b	:	IN STD_LOGIC := '0';
		byteena_a	:	IN STD_LOGIC_VECTOR(WIDTH_BYTEENA_A-1 DOWNTO 0) := (OTHERS => '1');
		byteena_b	:	IN STD_LOGIC_VECTOR(WIDTH_BYTEENA_B-1 DOWNTO 0) := (OTHERS => '1');
		clock0	:	IN STD_LOGIC := '1';
		clock1	:	IN STD_LOGIC := '1';
		clocken0	:	IN STD_LOGIC := '1';
		clocken1	:	IN STD_LOGIC := '1';
		clocken2	:	IN STD_LOGIC := '1';
		clocken3	:	IN STD_LOGIC := '1';
		data_a	:	IN STD_LOGIC_VECTOR(WIDTH_A-1 DOWNTO 0) := (OTHERS => '1');
		data_b	:	IN STD_LOGIC_VECTOR(WIDTH_B-1 DOWNTO 0) := (OTHERS => '1');
		eccstatus	:	OUT STD_LOGIC_VECTOR(2 DOWNTO 0);
		q_a	:	OUT STD_LOGIC_VECTOR(WIDTH_A-1 DOWNTO 0);
		q_b	:	OUT STD_LOGIC_VECTOR(WIDTH_B-1 DOWNTO 0);
		rden_a	:	IN STD_LOGIC := '1';
		rden_b	:	IN STD_LOGIC := '1';
		wren_a	:	IN STD_LOGIC := '0';
		wren_b	:	IN STD_LOGIC := '0'
	 ); 
	 END COMPONENT;
 BEGIN

	wire_w_lg_sclr4w(0) <= NOT sclr;
	wire_w_lg_sload_data31w(0) <= NOT sload_data;
	result <= ( result_wire(63 DOWNTO 0));
	result_valid <= dffe2a10;
	result_wire <= ( wire_accum7_result(35 DOWNTO 0) & wire_altshiftreg8_q(27 DOWNTO 0));
	sclr <= '0';
	wire_abs3_data <= ( wire_altshiftreg1_shiftout);
	wire_abs3_sign_bit <= wire_dffe5a_w_lg_q42w(0);
	wire_abs3_sload_data <= ( data_in(3 DOWNTO 0));
	abs3 :  memmult_abs_bla
	  PORT MAP ( 
		a_abs => dffe5a5,
		clock => clock,
		data => wire_abs3_data,
		result => wire_abs3_result,
		sign_bit => wire_abs3_sign_bit,
		sload => sload_data,
		sload_data => wire_abs3_sload_data
	  );
	wire_accum7_add_sub <= wire_dffe4a_w_lg_w_q_range54w55w(0);
	wire_dffe4a_w_lg_w_q_range54w55w(0) <= NOT dffe4a(3);
	wire_accum7_data <= ( wire_altsyncram6_q_a(35 DOWNTO 0));
	accum7 :  altaccumulate
	  GENERIC MAP (
		LPM_REPRESENTATION => "SIGNED",
		RIGHT_SHIFT_DISTANCE => 4,
		WIDTH_IN => 36,
		WIDTH_OUT => 37
	  )
	  PORT MAP ( 
		add_sub => wire_accum7_add_sub,
		clock => clock,
		data => wire_accum7_data,
		result => wire_accum7_result,
		sload => dffe2a2
	  );
	wire_altshiftreg1_data <= ( data_in(31 DOWNTO 4));
	altshiftreg1 :  memmult_altshiftreg_tda
	  PORT MAP ( 
		clock => clock,
		data => wire_altshiftreg1_data,
		load => sload_data,
		q => wire_altshiftreg1_q,
		shiftout => wire_altshiftreg1_shiftout
	  );
	altshiftreg8 :  memmult_altshiftreg_ji9
	  PORT MAP ( 
		clock => clock,
		q => wire_altshiftreg8_q,
		shiftin => wire_accum7_result(3 DOWNTO 0),
		shiftout => wire_altshiftreg8_shiftout
	  );
	altsyncram6 :  altsyncram
	  GENERIC MAP (
		INIT_FILE => "memmult.hex",
		OPERATION_MODE => "ROM",
		OUTDATA_REG_A => "CLOCK0",
		RAM_BLOCK_TYPE => "AUTO",
		WIDTH_A => 36,
		WIDTHAD_A => 4,
		INTENDED_DEVICE_FAMILY => "Cyclone"
	  )
	  PORT MAP ( 
		address_a => wire_abs3_result(3 DOWNTO 0),
		clock0 => clock,
		q_a => wire_altsyncram6_q_a
	  );
	PROCESS (clock)
	BEGIN
		IF (clock = '1' AND clock'event) THEN dffe2a0 <= (sload_data AND wire_w_lg_sclr4w(0));
		END IF;
	END PROCESS;
	PROCESS (clock)
	BEGIN
		IF (clock = '1' AND clock'event) THEN dffe2a1 <= (dffe2a0 AND wire_w_lg_sclr4w(0));
		END IF;
	END PROCESS;
	PROCESS (clock)
	BEGIN
		IF (clock = '1' AND clock'event) THEN dffe2a2 <= (dffe2a1 AND wire_w_lg_sclr4w(0));
		END IF;
	END PROCESS;
	wire_dffe2a_w_lg_q9w(0) <= NOT dffe2a2;
	PROCESS (clock)
	BEGIN
		IF (clock = '1' AND clock'event) THEN dffe2a3 <= (dffe2a2 AND wire_w_lg_sclr4w(0));
		END IF;
	END PROCESS;
	wire_dffe2a_w_lg_q10w(0) <= dffe2a3 AND wire_dffe2a_w_lg_q9w(0);
	PROCESS (clock)
	BEGIN
		IF (clock = '1' AND clock'event) THEN dffe2a4 <= (wire_dffe2a_w_lg_q10w(0) AND wire_w_lg_sclr4w(0));
		END IF;
	END PROCESS;
	wire_dffe2a_w_lg_q12w(0) <= dffe2a4 AND wire_dffe2a_w_lg_q9w(0);
	PROCESS (clock)
	BEGIN
		IF (clock = '1' AND clock'event) THEN dffe2a5 <= (wire_dffe2a_w_lg_q12w(0) AND wire_w_lg_sclr4w(0));
		END IF;
	END PROCESS;
	wire_dffe2a_w_lg_q14w(0) <= dffe2a5 AND wire_dffe2a_w_lg_q9w(0);
	PROCESS (clock)
	BEGIN
		IF (clock = '1' AND clock'event) THEN dffe2a6 <= (wire_dffe2a_w_lg_q14w(0) AND wire_w_lg_sclr4w(0));
		END IF;
	END PROCESS;
	wire_dffe2a_w_lg_q16w(0) <= dffe2a6 AND wire_dffe2a_w_lg_q9w(0);
	PROCESS (clock)
	BEGIN
		IF (clock = '1' AND clock'event) THEN dffe2a7 <= (wire_dffe2a_w_lg_q16w(0) AND wire_w_lg_sclr4w(0));
		END IF;
	END PROCESS;
	wire_dffe2a_w_lg_q18w(0) <= dffe2a7 AND wire_dffe2a_w_lg_q9w(0);
	PROCESS (clock)
	BEGIN
		IF (clock = '1' AND clock'event) THEN dffe2a8 <= (wire_dffe2a_w_lg_q18w(0) AND wire_w_lg_sclr4w(0));
		END IF;
	END PROCESS;
	wire_dffe2a_w_lg_q20w(0) <= dffe2a8 AND wire_dffe2a_w_lg_q9w(0);
	PROCESS (clock)
	BEGIN
		IF (clock = '1' AND clock'event) THEN dffe2a9 <= (wire_dffe2a_w_lg_q20w(0) AND wire_w_lg_sclr4w(0));
		END IF;
	END PROCESS;
	wire_dffe2a_w_lg_q22w(0) <= dffe2a9 AND wire_dffe2a_w_lg_q9w(0);
	PROCESS (clock)
	BEGIN
		IF (clock = '1' AND clock'event) THEN dffe2a10 <= (wire_dffe2a_w_lg_q22w(0) AND wire_w_lg_sclr4w(0));
		END IF;
	END PROCESS;
	PROCESS (clock)
	BEGIN
		IF (clock = '1' AND clock'event) THEN dffe4a <= ( dffe4a(2 DOWNTO 0) & wire_dffe5a_w_lg_q42w);
		END IF;
	END PROCESS;
	wire_dffe4a_w44w <= ( dffe4a(2 DOWNTO 0) & wire_dffe5a_w_lg_q42w);
	PROCESS (clock)
	BEGIN
		IF (clock = '1' AND clock'event) THEN dffe5a0 <= (data_in(31) AND sload_data);
		END IF;
	END PROCESS;
	wire_dffe5a_w_lg_q32w(0) <= dffe5a0 AND wire_w_lg_sclr4w(0);
	PROCESS (clock)
	BEGIN
		IF (clock = '1' AND clock'event) THEN dffe5a1 <= (wire_dffe5a_w_lg_q32w(0) AND wire_w_lg_sload_data31w(0));
		END IF;
	END PROCESS;
	wire_dffe5a_w_lg_q34w(0) <= dffe5a1 AND wire_w_lg_sclr4w(0);
	PROCESS (clock)
	BEGIN
		IF (clock = '1' AND clock'event) THEN dffe5a2 <= (wire_dffe5a_w_lg_q34w(0) AND wire_w_lg_sload_data31w(0));
		END IF;
	END PROCESS;
	wire_dffe5a_w_lg_q36w(0) <= dffe5a2 AND wire_w_lg_sclr4w(0);
	PROCESS (clock)
	BEGIN
		IF (clock = '1' AND clock'event) THEN dffe5a3 <= (wire_dffe5a_w_lg_q36w(0) AND wire_w_lg_sload_data31w(0));
		END IF;
	END PROCESS;
	wire_dffe5a_w_lg_q38w(0) <= dffe5a3 AND wire_w_lg_sclr4w(0);
	PROCESS (clock)
	BEGIN
		IF (clock = '1' AND clock'event) THEN dffe5a4 <= (wire_dffe5a_w_lg_q38w(0) AND wire_w_lg_sload_data31w(0));
		END IF;
	END PROCESS;
	wire_dffe5a_w_lg_q40w(0) <= dffe5a4 AND wire_w_lg_sclr4w(0);
	PROCESS (clock)
	BEGIN
		IF (clock = '1' AND clock'event) THEN dffe5a5 <= (wire_dffe5a_w_lg_q40w(0) AND wire_w_lg_sload_data31w(0));
		END IF;
	END PROCESS;
	wire_dffe5a_w_lg_q42w(0) <= dffe5a5 AND wire_w_lg_sload_data31w(0);

 END RTL; --memmult_altmemmult_v6q
--VALID FILE


LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY memmult IS
	PORT
	(
		clock		: IN STD_LOGIC ;
		data_in		: IN STD_LOGIC_VECTOR (31 DOWNTO 0);
		sload_data		: IN STD_LOGIC ;
		result		: OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
		result_valid		: OUT STD_LOGIC 
	);
END memmult;


ARCHITECTURE RTL OF memmult IS

	ATTRIBUTE synthesis_clearbox: boolean;
	ATTRIBUTE synthesis_clearbox OF RTL: ARCHITECTURE IS TRUE;
	SIGNAL sub_wire0	: STD_LOGIC ;
	SIGNAL sub_wire1	: STD_LOGIC_VECTOR (63 DOWNTO 0);



	COMPONENT memmult_altmemmult_v6q
	PORT (
			data_in	: IN STD_LOGIC_VECTOR (31 DOWNTO 0);
			clock	: IN STD_LOGIC ;
			result_valid	: OUT STD_LOGIC ;
			result	: OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
			sload_data	: IN STD_LOGIC 
	);
	END COMPONENT;

BEGIN
	result_valid    <= sub_wire0;
	result    <= sub_wire1(63 DOWNTO 0);

	memmult_altmemmult_v6q_component : memmult_altmemmult_v6q
	PORT MAP (
		data_in => data_in,
		clock => clock,
		sload_data => sload_data,
		result_valid => sub_wire0,
		result => sub_wire1
	);



END RTL;

-- ============================================================
-- CNX file retrieval info
-- ============================================================
-- Retrieval info: PRIVATE: COEFFICIENT0 STRING "1234"
-- Retrieval info: PRIVATE: COEFF_REPRESENTATION_COMBO STRING "SIGNED"
-- Retrieval info: PRIVATE: COUNT_C_COMBO STRING "32"
-- Retrieval info: PRIVATE: COUNT_D_COMBO STRING "32"
-- Retrieval info: PRIVATE: DATA_REPRESENTATION_COMBO STRING "SIGNED"
-- Retrieval info: PRIVATE: INTENDED_DEVICE_FAMILY STRING "Cyclone"
-- Retrieval info: PRIVATE: LOADABLE_COEFF STRING "0"
-- Retrieval info: PRIVATE: RAM_BLOCK_TYPE NUMERIC "0"
-- Retrieval info: PRIVATE: SCLR_CHECK STRING "0"
-- Retrieval info: PRIVATE: SYNTH_WRAPPER_GEN_POSTFIX STRING "0"
-- Retrieval info: PRIVATE: WIZMAN_OVERRIDE_CBX_GEN_MODE STRING "ON"
-- Retrieval info: CONSTANT: COEFFICIENT0 STRING "1234"
-- Retrieval info: CONSTANT: COEFF_REPRESENTATION STRING "SIGNED"
-- Retrieval info: CONSTANT: DATA_REPRESENTATION STRING "SIGNED"
-- Retrieval info: CONSTANT: INTENDED_DEVICE_FAMILY STRING "Cyclone"
-- Retrieval info: CONSTANT: MAX_CLOCK_CYCLES_PER_RESULT NUMERIC "8"
-- Retrieval info: CONSTANT: RAM_BLOCK_TYPE STRING "AUTO"
-- Retrieval info: CONSTANT: TOTAL_LATENCY NUMERIC "11"
-- Retrieval info: CONSTANT: WIDTH_C NUMERIC "32"
-- Retrieval info: CONSTANT: WIDTH_D NUMERIC "32"
-- Retrieval info: CONSTANT: WIDTH_R NUMERIC "64"
-- Retrieval info: USED_PORT: clock 0 0 0 0 INPUT NODEFVAL "clock"
-- Retrieval info: USED_PORT: data_in 0 0 32 0 INPUT NODEFVAL "data_in[31..0]"
-- Retrieval info: USED_PORT: result 0 0 64 0 OUTPUT NODEFVAL "result[63..0]"
-- Retrieval info: USED_PORT: result_valid 0 0 0 0 OUTPUT NODEFVAL "result_valid"
-- Retrieval info: USED_PORT: sload_data 0 0 0 0 INPUT NODEFVAL "sload_data"
-- Retrieval info: CONNECT: @data_in 0 0 32 0 data_in 0 0 32 0
-- Retrieval info: CONNECT: result_valid 0 0 0 0 @result_valid 0 0 0 0
-- Retrieval info: CONNECT: result 0 0 64 0 @result 0 0 64 0
-- Retrieval info: CONNECT: @sload_data 0 0 0 0 sload_data 0 0 0 0
-- Retrieval info: CONNECT: @clock 0 0 0 0 clock 0 0 0 0
-- Retrieval info: GEN_FILE: TYPE_NORMAL memmult.vhd TRUE FALSE
-- Retrieval info: GEN_FILE: TYPE_NORMAL memmult.inc FALSE FALSE
-- Retrieval info: GEN_FILE: TYPE_NORMAL memmult.cmp TRUE FALSE
-- Retrieval info: GEN_FILE: TYPE_NORMAL memmult.bsf TRUE FALSE
-- Retrieval info: GEN_FILE: TYPE_NORMAL memmult_inst.vhd FALSE FALSE
-- Retrieval info: LIB_FILE: altera_mf
-- Retrieval info: LIB_FILE: cyclone
